module ROM (
	input logic clk,
	input logic rst
);

endmodule
