module ROM (
	input logic clk,
	input logic rst,
	input logic [31:0] address,
	output logic [31:0] mem_out
);



endmodule
