module RAM (
	input logic clk,
	input logic rst
);

endmodule
