module ROM (
	input logic clk,
	input logic rst,
	input logic [31:0] PC,
	output logic [31:0] inst
);
	
	logic [31:0] instruction_set [0:407];
	
	initial begin
		instruction_set[0] = 32'hE3A08001;
		instruction_set[1] = 32'hE3A07003;
		instruction_set[2] = 32'hE3A09A02;
		instruction_set[3] = 32'hE3A0005A;
		instruction_set[4] = 32'hE5890008;
		instruction_set[5] = 32'hE3A0C000;
		instruction_set[6] = 32'hEB00001D;
		instruction_set[7] = 32'hEB000098;
		instruction_set[8] = 32'hEB000149;
		instruction_set[9] = 32'hEAFFFFFF;
		instruction_set[10] = 32'hEB0000C1;
		instruction_set[11] = 32'hEB000094;
		instruction_set[12] = 32'hE3580001;
		instruction_set[13] = 32'h0A000004;
		instruction_set[14] = 32'hE3580002;
		instruction_set[15] = 32'h0A000009;
		instruction_set[16] = 32'hE3580003;
		instruction_set[17] = 32'h0A00000E;
		instruction_set[18] = 32'hEAFFFFF6;
		instruction_set[19] = 32'hE357000A;
		instruction_set[20] = 32'hBAFFFFF4;
		instruction_set[21] = 32'hE3A08002;
		instruction_set[22] = 32'hEB000035;
		instruction_set[23] = 32'hEB00013A;
		instruction_set[24] = 32'hE3A07002;
		instruction_set[25] = 32'hEAFFFFEF;
		instruction_set[26] = 32'hE357000A;
		instruction_set[27] = 32'hBAFFFFED;
		instruction_set[28] = 32'hE3A08003;
		instruction_set[29] = 32'hEB000052;
		instruction_set[30] = 32'hEB000133;
		instruction_set[31] = 32'hE3A07002;
		instruction_set[32] = 32'hEAFFFFE8;
		instruction_set[33] = 32'hE357000A;
		instruction_set[34] = 32'hBAFFFFE6;
		instruction_set[35] = 32'hEB00016A;
		instruction_set[36] = 32'hEA000170;
		instruction_set[37] = 32'hE52DC004;
		instruction_set[38] = 32'hE3A0C064;
		instruction_set[39] = 32'hE3A00A01;
		instruction_set[40] = 32'hE3A02000;
		instruction_set[41] = 32'hE5802000;
		instruction_set[42] = 32'hE2800004;
		instruction_set[43] = 32'hE24CC001;
		instruction_set[44] = 32'hE35C0000;
		instruction_set[45] = 32'h1AFFFFFA;
		instruction_set[46] = 32'hE49DC004;
		instruction_set[47] = 32'hE3A00A01;
		instruction_set[48] = 32'hE3A03004;
		instruction_set[49] = 32'hE580307C;
		instruction_set[50] = 32'hE5803080;
		instruction_set[51] = 32'hE5803084;
		instruction_set[52] = 32'hE5803090;
		instruction_set[53] = 32'hE5803094;
		instruction_set[54] = 32'hE58030A8;
		instruction_set[55] = 32'hE58030B8;
		instruction_set[56] = 32'hE58030BC;
		instruction_set[57] = 32'hE58030C0;
		instruction_set[58] = 32'hE58030D0;
		instruction_set[59] = 32'hE58030E0;
		instruction_set[60] = 32'hE58030E4;
		instruction_set[61] = 32'hE58030E8;
		instruction_set[62] = 32'hE58030F8;
		instruction_set[63] = 32'hE5803108;
		instruction_set[64] = 32'hE580310C;
		instruction_set[65] = 32'hE3A03005;
		instruction_set[66] = 32'hE5803018;
		instruction_set[67] = 32'hE3A00C12;
		instruction_set[68] = 32'hE3A03008;
		instruction_set[69] = 32'hE5803000;
		instruction_set[70] = 32'hE3A03004;
		instruction_set[71] = 32'hE5803004;
		instruction_set[72] = 32'hE3A03000;
		instruction_set[73] = 32'hE5803008;
		instruction_set[74] = 32'hE3A030D7;
		instruction_set[75] = 32'hE580300C;
		instruction_set[76] = 32'hE12FFF1E;
		instruction_set[77] = 32'hE52DC004;
		instruction_set[78] = 32'hE3A0C064;
		instruction_set[79] = 32'hE3A00A01;
		instruction_set[80] = 32'hE3A02000;
		instruction_set[81] = 32'hE5802000;
		instruction_set[82] = 32'hE2800004;
		instruction_set[83] = 32'hE24CC001;
		instruction_set[84] = 32'h1AFFFFFB;
		instruction_set[85] = 32'hE49DC004;
		instruction_set[86] = 32'hE3A00A01;
		instruction_set[87] = 32'hE3A03004;
		instruction_set[88] = 32'hE5803000;
		instruction_set[89] = 32'hE580300C;
		instruction_set[90] = 32'hE5803018;
		instruction_set[91] = 32'hE5803024;
		instruction_set[92] = 32'hE5803058;
		instruction_set[93] = 32'hE580306C;
		instruction_set[94] = 32'hE5803078;
		instruction_set[95] = 32'hE5803084;
		instruction_set[96] = 32'hE5803090;
		instruction_set[97] = 32'hE580309C;
		instruction_set[98] = 32'hE58030F0;
		instruction_set[99] = 32'hE58030FC;
		instruction_set[100] = 32'hE5803108;
		instruction_set[101] = 32'hE5803114;
		instruction_set[102] = 32'hE5803120;
		instruction_set[103] = 32'hE5803134;
		instruction_set[104] = 32'hE5803168;
		instruction_set[105] = 32'hE5803174;
		instruction_set[106] = 32'hE5803180;
		instruction_set[107] = 32'hE580318C;
		instruction_set[108] = 32'hE3A03001;
		instruction_set[109] = 32'hE580302C;
		instruction_set[110] = 32'hE3A03002;
		instruction_set[111] = 32'hE5803030;
		instruction_set[112] = 32'hE12FFF1E;
		instruction_set[113] = 32'hE52DC004;
		instruction_set[114] = 32'hE3A0C064;
		instruction_set[115] = 32'hE3A01A01;
		instruction_set[116] = 32'hE3A02000;
		instruction_set[117] = 32'hE5812000;
		instruction_set[118] = 32'hE2811004;
		instruction_set[119] = 32'hE25CC001;
		instruction_set[120] = 32'h1AFFFFFB;
		instruction_set[121] = 32'hE49DC004;
		instruction_set[122] = 32'hE3A00A01;
		instruction_set[123] = 32'hE3A03004;
		instruction_set[124] = 32'hE5803000;
		instruction_set[125] = 32'hE5803004;
		instruction_set[126] = 32'hE5803020;
		instruction_set[127] = 32'hE5803024;
		instruction_set[128] = 32'hE5803028;
		instruction_set[129] = 32'hE5803040;
		instruction_set[130] = 32'hE580304C;
		instruction_set[131] = 32'hE580305C;
		instruction_set[132] = 32'hE5803060;
		instruction_set[133] = 32'hE5803064;
		instruction_set[134] = 32'hE5803068;
		instruction_set[135] = 32'hE5803084;
		instruction_set[136] = 32'hE58030A4;
		instruction_set[137] = 32'hE58030AC;
		instruction_set[138] = 32'hE58030C0;
		instruction_set[139] = 32'hE58030CC;
		instruction_set[140] = 32'hE58030E0;
		instruction_set[141] = 32'hE58030E8;
		instruction_set[142] = 32'hE5803108;
		instruction_set[143] = 32'hE5803124;
		instruction_set[144] = 32'hE5803128;
		instruction_set[145] = 32'hE580312C;
		instruction_set[146] = 32'hE5803130;
		instruction_set[147] = 32'hE5803140;
		instruction_set[148] = 32'hE580314C;
		instruction_set[149] = 32'hE5803164;
		instruction_set[150] = 32'hE5803168;
		instruction_set[151] = 32'hE580316C;
		instruction_set[152] = 32'hE5803188;
		instruction_set[153] = 32'hE580318C;
		instruction_set[154] = 32'hE3A03001;
		instruction_set[155] = 32'hE58130B4;
		instruction_set[156] = 32'hE3A03002;
		instruction_set[157] = 32'hE58130B0;
		instruction_set[158] = 32'hE12FFF1E;
		instruction_set[159] = 32'hE2877001;
		instruction_set[160] = 32'hE12FFF1E;
		instruction_set[161] = 32'hE52D0004;
		instruction_set[162] = 32'hE52D1004;
		instruction_set[163] = 32'hE52D2004;
		instruction_set[164] = 32'hE52D3004;
		instruction_set[165] = 32'hE52D4004;
		instruction_set[166] = 32'hE52DE004;
		instruction_set[167] = 32'hE3A00A01;
		instruction_set[168] = 32'hE3A01C12;
		instruction_set[169] = 32'hE3A02001;
		instruction_set[170] = 32'hE3A03004;
		instruction_set[171] = 32'hE0030793;
		instruction_set[172] = 32'hE3520000;
		instruction_set[173] = 32'h0A000009;
		instruction_set[174] = 32'hE7914003;
		instruction_set[175] = 32'hE3A050D7;
		instruction_set[176] = 32'hE1540005;
		instruction_set[177] = 32'h0A000005;
		instruction_set[178] = 32'hE0844000;
		instruction_set[179] = 32'hE3A05000;
		instruction_set[180] = 32'hE5845000;
		instruction_set[181] = 32'hE2833004;
		instruction_set[182] = 32'hE2422001;
		instruction_set[183] = 32'hEAFFFFF3;
		instruction_set[184] = 32'hE3A00A01;
		instruction_set[185] = 32'hE3A01C12;
		instruction_set[186] = 32'hE1A02007;
		instruction_set[187] = 32'hE3A03000;
		instruction_set[188] = 32'hE3A04001;
		instruction_set[189] = 32'hE3520000;
		instruction_set[190] = 32'h0A000006;
		instruction_set[191] = 32'hE7915003;
		instruction_set[192] = 32'hE0855000;
		instruction_set[193] = 32'hE5854000;
		instruction_set[194] = 32'hE3A04002;
		instruction_set[195] = 32'hE2833004;
		instruction_set[196] = 32'hE2422001;
		instruction_set[197] = 32'hEAFFFFF6;
		instruction_set[198] = 32'hE49DE004;
		instruction_set[199] = 32'hE49D4004;
		instruction_set[200] = 32'hE49D3004;
		instruction_set[201] = 32'hE49D2004;
		instruction_set[202] = 32'hE49D1004;
		instruction_set[203] = 32'hE49D0004;
		instruction_set[204] = 32'hE12FFF1E;
		instruction_set[205] = 32'hE52DE004;
		instruction_set[206] = 32'hEB00007B;
		instruction_set[207] = 32'hEB000022;
		instruction_set[208] = 32'hE3A06000;
		instruction_set[209] = 32'hE3A00C12;
		instruction_set[210] = 32'hE5901000;
		instruction_set[211] = 32'hEB00004B;
		instruction_set[212] = 32'hE3560000;
		instruction_set[213] = 32'hBA0000B9;
		instruction_set[214] = 32'hE3560F63;
		instruction_set[215] = 32'hCA0000B7;
		instruction_set[216] = 32'hE3A02A01;
		instruction_set[217] = 32'hE0823006;
		instruction_set[218] = 32'hE5934000;
		instruction_set[219] = 32'hE3540004;
		instruction_set[220] = 32'h0A0000B2;
		instruction_set[221] = 32'hE3540002;
		instruction_set[222] = 32'h0A0000B0;
		instruction_set[223] = 32'hE3540005;
		instruction_set[224] = 32'h0A00000A;
		instruction_set[225] = 32'hEB000003;
		instruction_set[226] = 32'hE3A00C12;
		instruction_set[227] = 32'hE5806000;
		instruction_set[228] = 32'hE49DE004;
		instruction_set[229] = 32'hE12FFF1E;
		instruction_set[230] = 32'hE3A00C12;
		instruction_set[231] = 32'hE1A01007;
		instruction_set[232] = 32'hE1A01101;
		instruction_set[233] = 32'hE0800001;
		instruction_set[234] = 32'hE1A02007;
		instruction_set[235] = 32'hEA000056;
		instruction_set[236] = 32'hEBFFFFB1;
		instruction_set[237] = 32'hEBFFFFF7;
		instruction_set[238] = 32'hE3A00C12;
		instruction_set[239] = 32'hE5806000;
		instruction_set[240] = 32'hEB000061;
		instruction_set[241] = 32'hE49DE004;
		instruction_set[242] = 32'hE12FFF1E;
		instruction_set[243] = 32'hE5994000;
		instruction_set[244] = 32'hE3A0204E;
		instruction_set[245] = 32'hE1540002;
		instruction_set[246] = 32'h0A000009;
		instruction_set[247] = 32'hE3A02020;
		instruction_set[248] = 32'hE1540002;
		instruction_set[249] = 32'h0A000006;
		instruction_set[250] = 32'hE3A0202D;
		instruction_set[251] = 32'hE1540002;
		instruction_set[252] = 32'h0A000003;
		instruction_set[253] = 32'hE3A02041;
		instruction_set[254] = 32'hE1540002;
		instruction_set[255] = 32'h0A000000;
		instruction_set[256] = 32'hE12FFF1E;
		instruction_set[257] = 32'hE5990000;
		instruction_set[258] = 32'hE5991004;
		instruction_set[259] = 32'hE3A0204E;
		instruction_set[260] = 32'hE1500002;
		instruction_set[261] = 32'h0A000009;
		instruction_set[262] = 32'hE3A02020;
		instruction_set[263] = 32'hE1500002;
		instruction_set[264] = 32'h0A000006;
		instruction_set[265] = 32'hE3A0202D;
		instruction_set[266] = 32'hE1500002;
		instruction_set[267] = 32'h0A00000A;
		instruction_set[268] = 32'hE3A02041;
		instruction_set[269] = 32'hE1500002;
		instruction_set[270] = 32'h0A000007;
		instruction_set[271] = 32'hEA00000E;
		instruction_set[272] = 32'hE3A0204E;
		instruction_set[273] = 32'hE1510002;
		instruction_set[274] = 32'h0A00000B;
		instruction_set[275] = 32'hE3A02020;
		instruction_set[276] = 32'hE1510002;
		instruction_set[277] = 32'h0A000008;
		instruction_set[278] = 32'hEA000006;
		instruction_set[279] = 32'hE3A0202D;
		instruction_set[280] = 32'hE1510002;
		instruction_set[281] = 32'h0A000004;
		instruction_set[282] = 32'hE3A02041;
		instruction_set[283] = 32'hE1510002;
		instruction_set[284] = 32'h0A000001;
		instruction_set[285] = 32'hEAFFFFFF;
		instruction_set[286] = 32'hE5890004;
		instruction_set[287] = 32'hE12FFF1E;
		instruction_set[288] = 32'hE5994004;
		instruction_set[289] = 32'hE3A0204E;
		instruction_set[290] = 32'hE1540002;
		instruction_set[291] = 32'h0A000016;
		instruction_set[292] = 32'hE3A02020;
		instruction_set[293] = 32'hE1540002;
		instruction_set[294] = 32'h0A000015;
		instruction_set[295] = 32'hE3A0202D;
		instruction_set[296] = 32'hE1540002;
		instruction_set[297] = 32'h0A000002;
		instruction_set[298] = 32'hE3A02041;
		instruction_set[299] = 32'hE1540002;
		instruction_set[300] = 32'h0A000006;
		instruction_set[301] = 32'hE1A02001;
		instruction_set[302] = 32'hE52DE004;
		instruction_set[303] = 32'hEB00004C;
		instruction_set[304] = 32'hE49DE004;
		instruction_set[305] = 32'hE3520000;
		instruction_set[306] = 32'h0A00005C;
		instruction_set[307] = 32'hEA00000A;
		instruction_set[308] = 32'hE1A02001;
		instruction_set[309] = 32'hE52DE004;
		instruction_set[310] = 32'hEB000045;
		instruction_set[311] = 32'hE49DE004;
		instruction_set[312] = 32'hE3520024;
		instruction_set[313] = 32'h0A000055;
		instruction_set[314] = 32'hEA000005;
		instruction_set[315] = 32'hE2416028;
		instruction_set[316] = 32'hE12FFF1E;
		instruction_set[317] = 32'hE2816028;
		instruction_set[318] = 32'hE12FFF1E;
		instruction_set[319] = 32'hE2416004;
		instruction_set[320] = 32'hE12FFF1E;
		instruction_set[321] = 32'hE2816004;
		instruction_set[322] = 32'hE12FFF1E;
		instruction_set[323] = 32'hE2400004;
		instruction_set[324] = 32'hE5903000;
		instruction_set[325] = 32'hE2804004;
		instruction_set[326] = 32'hE5843000;
		instruction_set[327] = 32'hE2422001;
		instruction_set[328] = 32'hE3520000;
		instruction_set[329] = 32'h1AFFFFF8;
		instruction_set[330] = 32'hE12FFF1E;
		instruction_set[331] = 32'hE3A00005;
		instruction_set[332] = 32'hE15C0000;
		instruction_set[333] = 32'h0A000003;
		instruction_set[334] = 32'hE3A00041;
		instruction_set[335] = 32'hE5890000;
		instruction_set[336] = 32'hE28CC001;
		instruction_set[337] = 32'hE12FFF1E;
		instruction_set[338] = 32'hE12FFF1E;
		instruction_set[339] = 32'hE52D1004;
		instruction_set[340] = 32'hE52D2004;
		instruction_set[341] = 32'hE52D3004;
		instruction_set[342] = 32'hE52D4004;
		instruction_set[343] = 32'hE52D5004;
		instruction_set[344] = 32'hE52D6004;
		instruction_set[345] = 32'hE52D7004;
		instruction_set[346] = 32'hE52DE004;
		instruction_set[347] = 32'hE52DC004;
		instruction_set[348] = 32'hE5992008;
		instruction_set[349] = 32'hE2822025;
		instruction_set[350] = 32'hE3A03049;
		instruction_set[351] = 32'hE0020392;
		instruction_set[352] = 32'hE20220FF;
		instruction_set[353] = 32'hE5892008;
		instruction_set[354] = 32'hE1A0A002;
		instruction_set[355] = 32'hEB00001E;
		instruction_set[356] = 32'hE2822061;
		instruction_set[357] = 32'hE1A0B002;
		instruction_set[358] = 32'hEB000021;
		instruction_set[359] = 32'hE3A03A01;
		instruction_set[360] = 32'hE3A0500A;
		instruction_set[361] = 32'hE004059A;
		instruction_set[362] = 32'hE084400B;
		instruction_set[363] = 32'hE3A05002;
		instruction_set[364] = 32'hE1A04514;
		instruction_set[365] = 32'hE0833004;
		instruction_set[366] = 32'hE5935000;
		instruction_set[367] = 32'hE3550000;
		instruction_set[368] = 32'h1AFFFFEA;
		instruction_set[369] = 32'hE3A05005;
		instruction_set[370] = 32'hE5835000;
		instruction_set[371] = 32'hE49DC004;
		instruction_set[372] = 32'hE49DE004;
		instruction_set[373] = 32'hE49D7004;
		instruction_set[374] = 32'hE49D6004;
		instruction_set[375] = 32'hE49D5004;
		instruction_set[376] = 32'hE49D4004;
		instruction_set[377] = 32'hE49D3004;
		instruction_set[378] = 32'hE49D2004;
		instruction_set[379] = 32'hE49D1004;
		instruction_set[380] = 32'hE12FFF1E;
		instruction_set[381] = 32'hE3A03028;
		instruction_set[382] = 32'hE1520003;
		instruction_set[383] = 32'hBA000001;
		instruction_set[384] = 32'hE0422003;
		instruction_set[385] = 32'hEAFFFFFB;
		instruction_set[386] = 32'hE12FFF1E;
		instruction_set[387] = 32'hE3A0C00A;
		instruction_set[388] = 32'hE15A000C;
		instruction_set[389] = 32'hBA000001;
		instruction_set[390] = 32'hE04AA00C;
		instruction_set[391] = 32'hEAFFFFFB;
		instruction_set[392] = 32'hE12FFF1E;
		instruction_set[393] = 32'hE3A0C00A;
		instruction_set[394] = 32'hE15B000C;
		instruction_set[395] = 32'hBA000001;
		instruction_set[396] = 32'hE04BB00C;
		instruction_set[397] = 32'hEAFFFFFB;
		instruction_set[398] = 32'hE12FFF1E;
		instruction_set[399] = 32'hEA000005;
		instruction_set[400] = 32'hE5901000;
		instruction_set[401] = 32'hE3A02A01;
		instruction_set[402] = 32'hE0823001;
		instruction_set[403] = 32'hE3A04008;
		instruction_set[404] = 32'hE5834000;
		instruction_set[405] = 32'hEAFFFFFF;
		instruction_set[406] = 32'hEAFFFFFE;
		instruction_set[407] = 32'h00000000;
	end
	
	always_ff @(posedge clk or posedge rst) begin
		if (rst)
			inst <= 32'h0;
		else if (PC >> 2 < 408)
			inst <= instruction_set[PC >> 2];
	end
	
endmodule
