module video_gen(
    input  logic [9:0] x,
    input  logic [9:0] y,
    input  logic blank_b,
    input  logic [3:0] matriz [9:0][9:0],
    output logic [7:0] r, g, b
);

    localparam CELL_SIZE   = 40;
    localparam GRID_WIDTH  = CELL_SIZE * 10;   // 400
    localparam GRID_HEIGHT = CELL_SIZE * 10;   // 400
    localparam SCREEN_WIDTH  = 640;
    localparam SCREEN_HEIGHT = 480;
    localparam OFFSET_X = (SCREEN_WIDTH - GRID_WIDTH) / 2;
    localparam OFFSET_Y = (SCREEN_HEIGHT - GRID_HEIGHT) / 2;

    logic [3:0] fila, col;
    logic [9:0] x_in_cell, y_in_cell;
    logic [3:0] valor;
    logic dentro_grid;

    assign dentro_grid = (x >= OFFSET_X && x < (OFFSET_X + GRID_WIDTH)) &&
                         (y >= OFFSET_Y && y < (OFFSET_Y + GRID_HEIGHT));

    assign col = (x - OFFSET_X) / CELL_SIZE;
    assign fila = (y - OFFSET_Y) / CELL_SIZE;
    assign x_in_cell = (x - OFFSET_X) % CELL_SIZE;
    assign y_in_cell = (y - OFFSET_Y) % CELL_SIZE;

    // Asignar valor de la celda de forma combinacional pura
    assign valor = (dentro_grid && blank_b) ? matriz[fila][col] : 4'd0;

    always_comb begin
        // Por defecto, pantalla negra
        r = 8'h00;
        g = 8'h00;
        b = 8'h00;

        if (blank_b && dentro_grid) begin
            if (x_in_cell == 0 || y_in_cell == 0) begin
                r = 8'h00; g = 8'h00; b = 8'h00; // bordes
            end else begin
                unique case (valor)
                    4'd0: begin r = 8'hFF; g = 8'hFF; b = 8'hFF; end // blanco
                    4'd1: begin r = 8'h00; g = 8'h80; b = 8'h00; end // verde oscuro
                    4'd2: begin r = 8'h90; g = 8'hEE; b = 8'h90; end // verde claro
                    4'd4: begin r = 8'h8B; g = 8'h45; b = 8'h13; end // café
                    4'd5: begin r = 8'hFF; g = 8'h00; b = 8'h00; end // rojo
						  4'd8: begin r = 8'hFF; g = 8'hFF; b = 8'h00; end // rojo
                    default: begin r = 8'hC0; g = 8'hC0; b = 8'hC0; end // gris claro
                endcase
            end
        end
    end

endmodule
