module ControlUnit (
	
);

	
endmodule
